PROBLEMA 1.3
V1 4 0 AC 40 45
V2 4 3 AC 80 45
R1 0 1 20
R2 1 5 10
R3 3 2 20
L 4 5 31.83m
C 2 1 79.57u
.AC LIN 1 50 50
.PRINT AC I(V1) IP(V1) I(V2) IP(V2) I(R1) IP(R1) I(R2) IP(R2) I(R3) IP(R3) I(L) IP(L) I(C) IP(C)
.END

; p este phase
; .PROBE -> pentru editor grafic