CIRCUIT T PODIT
* acesta este ;primul circuit simulat
VPOLARIZARE 1 0 12
* ce a fost mai sus este sursa de tensiune intre nodurile 1 si 0 si are 12 V
R1 1 2 10 
* rezistenmta 1 se afla intre nodurile 1 si 2 si arte 10 ohmi
* asemanator e si la restul =)
R2 2 0 10
R3 2 3 5
R4 1 3 5
* .OP este pentru aflarea valorii potentialelor
* .END este pentru final de fisier
.OP
.END


