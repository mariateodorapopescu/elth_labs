TEMA 3
V1 3 4 90
V2 5 4 90
V3 1 4 50
I1 2 1 5
R1 3 0 10
R2 1 0 5
R3 5 0 10
R4 2 3 30
R5 2 4 10
.op
.dc V3 50 50 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) V(I1) I(V3)
.end
