TEMA 2
V1 5 1 50
V2 3 2 30
V3 5 4 90
I1 1 0 2
R1 0 4 25
R2 5 2 12
R3 1 2 10
R4 4 3 10
R5 0 5 10
.op
.dc V1 50 50 1
.print dc I(R1) I(R2) I(R3) I(R4) I(R5) I(V1) I(V2) I(V3) V(I1)
.end
