EXERCITIUL_A
*
R1 1 0 2
R2 0 4 1
R3 0 5 4
R5 2 3 2
*
V1 1 2 12
V3 3 5 4
I4 0 2 4
H2 4 3 V1 -2
*
.dc V1 12 12 1
.print dc I(R1) I(R2) I(R3) I(R5) V(I4)
.op
*
.end
