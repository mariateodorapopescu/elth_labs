PROBLEMA 3.1
Vin 1 0 AC 1
R 1 2 100
L 2 3 25.33m
C 3 0 1u
.AC lin 1000 100Hz 10kHz
.PROBE
.END