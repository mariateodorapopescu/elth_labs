EXERCITIUL_C
*
R1 0 1 2
R2 2 3 2 
R3 1 3 2
R4 4 3 2
* 
V1 4 0 12
V2 1 2 6
*
G5 4 3 1 0 1
*
.dc V1 12 12 1
.print dc I(R1) I(R2) I(R3) I(R4) V(G5)
.op
*
.end

